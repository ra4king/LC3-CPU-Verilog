library verilog;
use verilog.vl_types.all;
entity LC3_CPU_Test is
end LC3_CPU_Test;
